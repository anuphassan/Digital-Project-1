module de10_test(
output f,
input a,
input b
);
and(f, a, b); // f = ab
endmodule